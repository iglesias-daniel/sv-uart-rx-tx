module top (

);



endmodule

