module uart_rx #(

) (

);



endmodule